// Copyright Antmicro 2023
// SPDX-License-Identifier: Apache-2.0

module phy
  import top_pkg::*;
  import tlul_pkg::*;
(
    input  wire        clk,
    input  wire        rst,
    output wire        clk_idelay,
    output wire        rst_idelay,
    output wire        clk_sys,
    output wire        rst_sys,
    output wire        clk_sys2x,
    output wire        rst_sys2x,
    output wire        clk_sys8x,
    output wire        rst_sys8x,

    output wire [ 5:0] ddram_ca,
    output wire        ddram_cs,
    inout  wire [15:0] ddram_dq,
    inout  wire [ 1:0] ddram_dqs_p,
    inout  wire [ 1:0] ddram_dqs_n,
    inout  wire [ 1:0] ddram_dmi,
    output wire        ddram_clk_p,
    output wire        ddram_clk_n,
    output wire        ddram_cke,
    output wire        ddram_odt,
    output wire        ddram_reset_n,
    input  wire        dfi_cke_p0,
    input  wire        dfi_reset_n_p0,
    input  wire        dfi_mode_2n_p0,
    output wire        dfi_alert_n_w0,
    input  wire [16:0] dfi_address_p0,
    input  wire [ 5:0] dfi_bank_p0,
    input  wire        dfi_cas_n_p0,
    input  wire        dfi_cs_n_p0,
    input  wire        dfi_ras_n_p0,
    input  wire        dfi_act_n_p0,
    input  wire        dfi_odt_p0,
    input  wire        dfi_we_n_p0,
    input  wire [31:0] dfi_wrdata_p0,
    input  wire        dfi_wrdata_en_p0,
    input  wire [ 3:0] dfi_wrdata_mask_p0,
    input  wire        dfi_rddata_en_p0,
    output wire [31:0] dfi_rddata_w0,
    output wire        dfi_rddata_valid_w0,
    input  wire        dfi_cke_p1,
    input  wire        dfi_reset_n_p1,
    input  wire        dfi_mode_2n_p1,
    output wire        dfi_alert_n_w1,
    input  wire [16:0] dfi_address_p1,
    input  wire [ 5:0] dfi_bank_p1,
    input  wire        dfi_cas_n_p1,
    input  wire        dfi_cs_n_p1,
    input  wire        dfi_ras_n_p1,
    input  wire        dfi_act_n_p1,
    input  wire        dfi_odt_p1,
    input  wire        dfi_we_n_p1,
    input  wire [31:0] dfi_wrdata_p1,
    input  wire        dfi_wrdata_en_p1,
    input  wire [ 3:0] dfi_wrdata_mask_p1,
    input  wire        dfi_rddata_en_p1,
    output wire [31:0] dfi_rddata_w1,
    output wire        dfi_rddata_valid_w1,
    input  wire        dfi_cke_p2,
    input  wire        dfi_reset_n_p2,
    input  wire        dfi_mode_2n_p2,
    output wire        dfi_alert_n_w2,
    input  wire [16:0] dfi_address_p2,
    input  wire [ 5:0] dfi_bank_p2,
    input  wire        dfi_cas_n_p2,
    input  wire        dfi_cs_n_p2,
    input  wire        dfi_ras_n_p2,
    input  wire        dfi_act_n_p2,
    input  wire        dfi_odt_p2,
    input  wire        dfi_we_n_p2,
    input  wire [31:0] dfi_wrdata_p2,
    input  wire        dfi_wrdata_en_p2,
    input  wire [ 3:0] dfi_wrdata_mask_p2,
    input  wire        dfi_rddata_en_p2,
    output wire [31:0] dfi_rddata_w2,
    output wire        dfi_rddata_valid_w2,
    input  wire        dfi_cke_p3,
    input  wire        dfi_reset_n_p3,
    input  wire        dfi_mode_2n_p3,
    output wire        dfi_alert_n_w3,
    input  wire [16:0] dfi_address_p3,
    input  wire [ 5:0] dfi_bank_p3,
    input  wire        dfi_cas_n_p3,
    input  wire        dfi_cs_n_p3,
    input  wire        dfi_ras_n_p3,
    input  wire        dfi_act_n_p3,
    input  wire        dfi_odt_p3,
    input  wire        dfi_we_n_p3,
    input  wire [31:0] dfi_wrdata_p3,
    input  wire        dfi_wrdata_en_p3,
    input  wire [ 3:0] dfi_wrdata_mask_p3,
    input  wire        dfi_rddata_en_p3,
    output wire [31:0] dfi_rddata_w3,
    output wire        dfi_rddata_valid_w3,
    input  wire        dfi_cke_p4,
    input  wire        dfi_reset_n_p4,
    input  wire        dfi_mode_2n_p4,
    output wire        dfi_alert_n_w4,
    input  wire [16:0] dfi_address_p4,
    input  wire [ 5:0] dfi_bank_p4,
    input  wire        dfi_cas_n_p4,
    input  wire        dfi_cs_n_p4,
    input  wire        dfi_ras_n_p4,
    input  wire        dfi_act_n_p4,
    input  wire        dfi_odt_p4,
    input  wire        dfi_we_n_p4,
    input  wire [31:0] dfi_wrdata_p4,
    input  wire        dfi_wrdata_en_p4,
    input  wire [ 3:0] dfi_wrdata_mask_p4,
    input  wire        dfi_rddata_en_p4,
    output wire [31:0] dfi_rddata_w4,
    output wire        dfi_rddata_valid_w4,
    input  wire        dfi_cke_p5,
    input  wire        dfi_reset_n_p5,
    input  wire        dfi_mode_2n_p5,
    output wire        dfi_alert_n_w5,
    input  wire [16:0] dfi_address_p5,
    input  wire [ 5:0] dfi_bank_p5,
    input  wire        dfi_cas_n_p5,
    input  wire        dfi_cs_n_p5,
    input  wire        dfi_ras_n_p5,
    input  wire        dfi_act_n_p5,
    input  wire        dfi_odt_p5,
    input  wire        dfi_we_n_p5,
    input  wire [31:0] dfi_wrdata_p5,
    input  wire        dfi_wrdata_en_p5,
    input  wire [ 3:0] dfi_wrdata_mask_p5,
    input  wire        dfi_rddata_en_p5,
    output wire [31:0] dfi_rddata_w5,
    output wire        dfi_rddata_valid_w5,
    input  wire        dfi_cke_p6,
    input  wire        dfi_reset_n_p6,
    input  wire        dfi_mode_2n_p6,
    output wire        dfi_alert_n_w6,
    input  wire [16:0] dfi_address_p6,
    input  wire [ 5:0] dfi_bank_p6,
    input  wire        dfi_cas_n_p6,
    input  wire        dfi_cs_n_p6,
    input  wire        dfi_ras_n_p6,
    input  wire        dfi_act_n_p6,
    input  wire        dfi_odt_p6,
    input  wire        dfi_we_n_p6,
    input  wire [31:0] dfi_wrdata_p6,
    input  wire        dfi_wrdata_en_p6,
    input  wire [ 3:0] dfi_wrdata_mask_p6,
    input  wire        dfi_rddata_en_p6,
    output wire [31:0] dfi_rddata_w6,
    output wire        dfi_rddata_valid_w6,
    input  wire        dfi_cke_p7,
    input  wire        dfi_reset_n_p7,
    input  wire        dfi_mode_2n_p7,
    output wire        dfi_alert_n_w7,
    input  wire [16:0] dfi_address_p7,
    input  wire [ 5:0] dfi_bank_p7,
    input  wire        dfi_cas_n_p7,
    input  wire        dfi_cs_n_p7,
    input  wire        dfi_ras_n_p7,
    input  wire        dfi_act_n_p7,
    input  wire        dfi_odt_p7,
    input  wire        dfi_we_n_p7,
    input  wire [31:0] dfi_wrdata_p7,
    input  wire        dfi_wrdata_en_p7,
    input  wire [ 3:0] dfi_wrdata_mask_p7,
    input  wire        dfi_rddata_en_p7,
    output wire [31:0] dfi_rddata_w7,
    output wire        dfi_rddata_valid_w7,

    input  tlul_pkg::tl_h2d_t tl_i,
    output tlul_pkg::tl_d2h_t tl_o
);

  wire [ 9:0] csr_adr;
  wire        csr_we;
  wire [31:0] csr_dat_w;
  wire [31:0] csr_dat_r;

  phy_core u_phy_core (.*);

  tlul_adapter_reg #(
      .RegAw(top_pkg::TL_AW),
      .RegDw(top_pkg::TL_DW)
  ) u_tlul_adapter_reg (
      .clk_i (clk),
      .rst_ni(~rst),

      .tl_i(tl_i),
      .tl_o(tl_o),

      .en_ifetch_i (MuBi4True),
      .intg_error_o(), // unused

      .re_o(), // unused
      .we_o(csr_we),
      .addr_o(csr_adr),
      .wdata_o(csr_dat_w),
      .be_o({top_pkg::TL_DBW{1'b1}}),
      .busy_i(1'b0),
      .rdata_i(csr_dat_r),
      .error_i(1'b0)
  );

endmodule
